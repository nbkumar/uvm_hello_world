package my_package;
	import uvm_pkg::*;

	class env extends uvm_env;
	endclass

	class test extends uvm_test;
	endclass
endpackage 
